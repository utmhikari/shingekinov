module main

import shingeki

fn main() {
	mut server := shingeki.server()
	server.start()
}